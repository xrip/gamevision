� ����L `� ���  � ��� `�@�  6��@�  2�`��,� � � �� � �?� � ��� � � �� � �?� `  � l�� � �� �� � � %��L|�L
�� �� 6��� �  �� ��� �  R��� �L��� �� Ɇ�  R��� �  6���� �� 6��@�  �� 6��� �  6�� �0 �� �� 6��	� �  �� �� 6�� ���  [��� �q � Li� �`  � V�� � � � � � �  6�� �� ��L5�L��� �� 6��� �  ���  �  ��� �  6��� �  ���   ���   ��� � �  M� �� ��i ��i�� 6���  [� ��� � � H� � hL� �`  ��� �  6�� � �� 6��� �  �� F� 6�� �8 �� �� 6���� �� 6�� � 6��  ���   ���  � ؇`  ��� �  6�� � ���   �� � � � ���   ��� �   � ��� �  6�� � � ܉�LT�� � ��� � � � � � �  6��� �  ��Lt�Lǂ� � �  6��� �  w���   ���   ���   ��� �  6��� �  }��  �� ��� � � H� � hLZ� ݇` _� ��ީ � � � �� � �� � ��� L��� � � � � � ��� � �	 �A���
 � � �؍ � ��� �ͩ�� �	 �O� �
 � � �؍ � ��� � �' � )��L��� �   6���  ���  燠 � � �% �� �ީ � � � �� � ��� L� ʇ`�  ��   �� � �� �� F� 6�� � ���   �� � � 6�� � 쉢   � V� � ���   ���  �L��� �   Ɇ� )��L��� � � %��L�� � �L�� ��L���� �  6��� �  F� }��LS��� �  6��� �  }��L\�� � �L`�� ��Lh�L����   ���   ��  ���� � H�� h��   ���   �� �� *�L��� �   Ɇ� )���L��� �   Ɇ� )��L݄�� � �� � *�L愢 � �Lꄢ ��L=���   ���   ��  ���� � H:�� h��   ���   �� �� *�L(�� �   Ɇ� )���L��� �   Ɇ� )��Lb��� � �  ��Lk�� � �Lo�� ��L���� � H:�� h� ��� ��   ���  � *�L��� �   Ɇ� )���L��� �   Ɇ� )��Lᅠ� �  6��� �  F� ��Lꅢ � �L ��L1��� � H�� h� ��� ��   ���  � *�L�� �   Ɇ� )���L��� �   Ɇ� )���L���� �  6�� � �� 6��� �  ���   �� � �  6���  ���  燠�  ˂ ��L� ݇`� r �� ���r �� ���`�H�e � ��h`�
&�`�
&
&
&�`I�H�I��h`� ����L `�����	� �
���ک��� ����
����	������` �� ކ� � � �  � �� ҆L"�H�' )��$ �&�' )��% �%h@�'@8���`�8���`� ��� `� 8�� �`�`� 8�� �`�`� �  ��L�� ��� � �� ��� � ��8��	��i�	`P�I�	`��e��`� ��`�� �� � �� �`� �`�L���L���L����	� �`���	����`�� ��� `�� �`��� �`��0�� �`�� �`��� �`�ۢ �*`��� ��� Ç��� �	�� �Ff�	�����	�e�
�	e������
ȑ�
����	��������
��LÇ���.� ���	�'��Ff�e��	e��fjff����`Lֈ�	�����L��� ����	��F�e��	e��fjf��몥`F�ejf�����`�� �	�� �Lʇ� � � �� � � `�� � `� � H� 8�� ����� h�� `� �`� � �H�� h`�H�� �	� ��Ȋ��h�Lʇ� 8I�r �H�I�q �hL��� �� � ����	`� ����&	*&��������������`&	*��������`� �  ��L+��  ��L%�� �� � ����`�%���	� �� �
�����	���������`                  < <        6 6             6 6  6  6 6    >   0       c 3   f c    6  n ; 3 n                                    f < � < f         ?                          ?                       ` 0        > c s { o g >         ?    3 0   3 ?    3 0  0 3    8 < 6 3  0 x   ?   0 0 3        3 3    ? 3 0        3 3  3 3     3 3 > 0                                         ?     ?        0       3 0        > c { { {       3 3 ? 3 3   ? f f > f f ?   < f    f <    6 f f f 6     F    F     F        < f   s f |   3 3 3 ? 3 3 3            x 0 0 0 3 3    g f 6  6 f g       F f    c w   k c c   c g o { s c c    6 c c c 6    ? f f >       3 3 3 ;  8   ? f f > 6 f g    3   8 3    ? -        3 3 3 3 3 3 ?   3 3 3 3 3     c c c k  w c   c c 6   6 c   3 3 3        c 1  L f                 0 ` @              6 c                       �                   0 > 3 n      > f f ;        3  3    8 0 0 > 3 3 n        3 ?      6            n 3 3 > 0    6 n f f g             0   0 0 0 3 3    f 6  6 g                3   k c        3 3 3 3        3 3 3        ; f f >       n 3 3 > 0 x     ; n f         >   0      >   ,        3 3 3 3 n       3 3 3         c k   6       c 6  6 c       3 3 3 > 0      ?   & ?   8      8                8      n ;                            ���������������! ������`������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ɍ& L���B���%�